// Interface
interface intf();
  logic a;
  logic b;
  logic c_in;
  logic sum;
  logic c_out;
  endinterface
