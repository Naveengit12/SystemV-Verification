// interface code

interface intf;
  logic clk;
  logic rstn;
  logic up_down;
  logic [2:0]count;
endinterface
