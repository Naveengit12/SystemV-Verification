// interface

interface intf(input clk, rstn);
//   logic clk;
//   logic rstn;
  logic d;
  logic q;
  logic q_;
endinterface
